library verilog;
use verilog.vl_types.all;
entity CODE6B_vlg_sample_tst is
    port(
        clk_in          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end CODE6B_vlg_sample_tst;
