library verilog;
use verilog.vl_types.all;
entity CODE6B_vlg_vec_tst is
end CODE6B_vlg_vec_tst;
